module block_rom ( input [7:0]	addr,
						output [15:0]	data
					 );

    parameter ADDR_WIDTH = 11;
    parameter DATA_WIDTH = 16;
    parameter BLOCKS_NUM = 2;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0: (16*BLOCKS_NUM - 1)][DATA_WIDTH-1:0] BLOCK_ROM = 
    {
        // code 0x0
        16'b1111111111111111, // 0
        16'b1111111111111111, // 1
        16'b1111111111111111, // 2
        16'b1111111111111111, // 5
        16'b1111111111111111, // 4
        16'b1111111111111111, // 6
        16'b1111111111111111, // 3
        16'b1111111111111111, // 7      // Block
        16'b1111111111111111, // 8
        16'b1111111111111111, // 9
        16'b1111111111111111, // a
        16'b1111111111111111, // b
        16'b1111111111111111, // c
        16'b1111111111111111, // d
        16'b1111111111111111, // e
        16'b1111111111111111, // f

        // code 0x1
        16'b0000000000000000, // 0
        16'b0000000000000000, // 1
        16'b0000000000000000, // 2
        16'b0000000000000000, // 5
        16'b0000000000000000, // 4
        16'b0000000000000000, // 6
        16'b0000000000000000, // 3
        16'b0000000000000000, // 7      // Background
        16'b0000000000000000, // 8
        16'b0000000000000000, // 9
        16'b0000000000000000, // a
        16'b0000000000000000, // b
        16'b0000000000000000, // c
        16'b0000000000000000, // d
        16'b0000000000000000, // e
        16'b0000000000000000 // f

        // code 0x2
        
        };

	assign data = BLOCK_ROM[addr];

endmodule  